OTA Integrator
VP 7 0 DC 12V
VN 4 0 DC -12V
VIN 2 0 PULSE(2 -2 0 1NS 1NS 0.05S 0.1S)
IB 5 0 DC 1uA
X 0 2 6 7 4 5 OTA1
C1 6 0 0.001UF
.LIB C:\Cadence\SPB_16.6\tools\pspice\OTA1.LIB
.TRAN 1MS 1V
.PROBE
.END