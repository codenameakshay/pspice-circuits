*Notch Filter
R0 1 2 10K
R1 1 3 10K
R2 2 6 20K
R3 5 10 10K
R4 10 0 10K
C1 3 5 10NF
C2 8 10 10NF
VP 7 0 15V
VN 4 0 -15V
X1 3 2 7 4 6 UA741
X2 5 8 7 4 8 UA741
VIN 1 0 AC 1MV
.LIB NOM.LIB
.AC DEC 100 1 100K
.PROBE
.END