AC ANALYSIS
R1 4 3 2K
R2 3 0 2K
R3 3 6 2K
R4 7 9 0.5K
R5 9 6 0.5K
R6 2 0 2K
R7 2 6 0.5K
X1 1 2 4 OPAMP1
X2 1 3 7 OPAMP1
X3 1 9 6 OPAMP1
.LIB C:\Cadence\SPB_16.6\tools\pspice\OPAMP1.LIB
VIN 1 0 AC 0.1V
.AC DEC 50 1 1MEG
.PROBE
.END