Simple Current Mirror
Q1 2 2 0 Q2N2222
Q2 3 2 0 Q2N2222
R0 1 2 9.3K
*VCC 1 0 DC 10V
V0 3 0 DC 2V
.PROBE
.LIB NOM.LIB
IIN 1 0 DC 1UA
.DC LIN IIN 1UA 1MA 1UA
*.DC LIN V0 1 2 0.1
.END