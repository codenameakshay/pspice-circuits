*Log-AntiLog Circuit
R1 1 2 1K
R2 10 9 1K
R3 5 4 1K
R4 7 13 1K
Q1 2 0 3 Q2N2222
Q2 7 8 6 Q2N2222
Q3 4 3 6 Q2N2222
Q4 9 0 8 Q2N2222
X1 0 2 11 12 3 UA741
X2 0 4 11 12 6 UA741
X3 0 9 11 12 8 UA741
X4 0 7 11 12 13 UA741
V1 1 0 1V
V2 10 0 1V
V3 5 0 1V
VDD 11 0 15V
VSS 12 0 -15V
.DC V2 -10 10 0.01V
.PROBE
.LIB NOM.LIB
.END
