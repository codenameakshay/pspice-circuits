Integrator
R1 1 2 2.5K
C1 2 6 10U
VIN 1 0 PULSE(2 -2 0 1NS 1NS 0.05S 0.1S)
VP 7 0 DC 12V
VN 4 0 DC -12V
X 0 2 7 4 6 UA741
.LIB NOM.LIB
.TRAN 1MS 1S
.PROBE
.END