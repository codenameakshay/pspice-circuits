*COMPENSATED INVERTING AMPLIFIER *
X1 0 3 4 5 6 UA741
X2 6 3 7 8 9 UA741
R1 1 3 1000
R2 3 9 1000
V1 4 0 DC 12V
V2 0 5 DC 12V
V3 7 0 DC 12V
V4 0 8 DC 12V
VIN 1 0 AC 100MV
.LIB NOM.LIB
.AC DEC 20 1HZ 100MEG
.PROBE
.END