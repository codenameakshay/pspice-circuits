*COMPENSATED INVERTING AMPLIFIER 2 *
X1 0 2 3 4 5 UA741
X2 5 6 7 8 9 UA741
R1 5 6 10K
R2 6 9 10K
R3 9 2 10K
R4 1 2 10K
VIN 1 0 AC 100MV
V1 3 0 DC 12V
V2 0 4 DC 12V
V3 7 0 DC 12V
V4 0 8 DC 12V
.LIB NOM.LIB
.AC DEC 20 1HZ 100MEG
.PROBE
.END