*INVERTING AMPLIFIER *
X1 0 2 3 4 5 UA741
R1 1 2 1000
R2 2 5 1000
V1 3 0 DC 12
V2 0 4 DC 12
VIN 1 0 AC 100MV
.AC DEC 20 1HZ 100MEG
.LIB NOM.LIB
.PROBE
.END