Differentiator
R1 2 6 0.5K
C1 1 2 10U
VIN 1 0 PWL(0 0 0.5MS 5 1MS 0 1.5MS 5 2MS 0 2.5MS 5 3MS 0 3.5MS 5 4MS 0)
VP 7 0 DC 12V
VN 4 0 DC -12V
X 0 2 7 4 6 UA741
.LIB NOM.LIB
.TRAN 10NS 4MS
.PROBE
.END